* /home/drako/applications/eSim-2.1/library/SubcircuitLibrary/and_gate/and_gate.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Jun 29 15:22:30 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M2  Net-_M1-Pad3_ Net-_M1-Pad2_ Net-_M2-Pad3_ Net-_M2-Pad3_ mosfet_n		
M3  Net-_M2-Pad3_ Net-_M3-Pad2_ GND GND mosfet_n		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad1_ mosfet_p		
M4  Net-_M1-Pad1_ Net-_M3-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad1_ mosfet_p		
M5  Net-_M5-Pad1_ Net-_M1-Pad3_ GND GND mosfet_n		
M6  Net-_M1-Pad1_ Net-_M1-Pad3_ Net-_M5-Pad1_ Net-_M1-Pad1_ mosfet_p		
U1  Net-_M1-Pad2_ Net-_M3-Pad2_ Net-_M5-Pad1_ PORT		
v1  Net-_M1-Pad1_ GND 3.3v		

.end
