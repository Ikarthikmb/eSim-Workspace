* /home/drako/eSim-Workspace/wstage2/wstage2.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Jun 29 23:26:11 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
x3  /r0 /p0 Net-_x3-Pad3_ and_gate		
U1  /q1 /q0 /q2 /q3 /p1 /p2 /p0 /p3 /r0 /s4 /s0 /s1 /s2 /s3 PORT		
x5  Net-_x3-Pad3_ /q0 /s0 Net-_x5-Pad4_ halfadder		
x2  /r0 /p2 Net-_x2-Pad3_ and_gate		
x4  /r0 /p3 Net-_x4-Pad3_ and_gate		
x1  /r0 /p1 Net-_x1-Pad3_ and_gate		
x6  Net-_x1-Pad3_ /q1 Net-_x5-Pad4_ /s1 Net-_x6-Pad5_ fulladder		
x7  Net-_x2-Pad3_ /q2 Net-_x6-Pad5_ /s2 Net-_x7-Pad5_ fulladder		
x8  Net-_x4-Pad3_ /q3 Net-_x7-Pad5_ /s3 /s4 fulladder		

.end
