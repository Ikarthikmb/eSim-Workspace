* /home/drako/esim-workspace/wallace2tree/wallace2tree.cir

.include halfadder.sub
.include and_gate.sub
x1 b0 a0 z0 halfadder
x2 b0 a1 net-_x2-pad3_ halfadder
x3 b1 a0 net-_x3-pad3_ and_gate
x1 net-_x3-pad3_ net-_x2-pad3_ z1 net-_x1-pad4_ halfadder
x4 b1 a1 net-_x4-pad3_ and_gate
x2 net-_x1-pad4_ net-_x4-pad3_ z2 z3 halfadder
* u1  a0 a1 b0 b1 z0 z1 z2 z3 port

v2 a_in gnd pulse 0 1.8 0 0.1n 0.1n 5n 10n 
v3 b_in gnd pulse 0 1.8 0 0.1n 0.1n 10n 20n 
v4 a_in gnd pulse 0 1.8 0 0.1n 0.1n 20n 40n 
v5 b_in gnd pulse 0 1.8 0 0.1n 0.1n 40n 80n 

.tran 0.1n 80n

* Control Statements 
.control
run
plot z0 z1 z2 z3
print allv > plot_data_v.txt
print alli > plot_data_i.txt
.endc
.end
