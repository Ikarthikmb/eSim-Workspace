* /home/drako/applications/eSim-2.1/library/SubcircuitLibrary/wallace2tree/wallace2tree.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed Jun 30 01:29:03 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
x2  /b0 /a0 /z0 and_gate		
x1  /b0 /a1 Net-_x1-Pad3_ and_gate		
x3  /b1 /a0 Net-_x3-Pad3_ and_gate		
x4  /b1 /a1 Net-_x4-Pad3_ and_gate		
x5  Net-_x3-Pad3_ Net-_x1-Pad3_ /z1 Net-_x5-Pad4_ halfadder		
x6  Net-_x5-Pad4_ Net-_x4-Pad3_ /z2 /z3 halfadder		
U1  /a1 /a0 /b0 /b1 /z0 /z1 /z2 /z3 PORT		

.end
