AND GATE

* /home/drako/eSim-Workspace/prelayout/and_gate.cir

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

xm2  net-_m1-pad3_ a_in net-_m2-pad3_ net-_m2-pad3_ sky130_fd_pr__nfet_01v8 w=1 l=0.5
xm3  net-_m2-pad3_ b_in gnd gnd sky130_fd_pr__nfet_01v8 w=1 l=0.5
xm5  and_out net-_m1-pad3_ gnd gnd sky130_fd_pr__nfet_01v8 w=1 l=0.5
xm1  vcc a_in net-_m1-pad3_ vcc sky130_fd_pr__pfet_01v8 w=1 l=0.5
xm4  vcc b_in net-_m1-pad3_ vcc sky130_fd_pr__pfet_01v8 w=1 l=0.5
xm6  vcc vcc and_out and_out sky130_fd_pr__pfet_01v8 w=1 l=0.5

v3 vcc gnd dc 3.3
v1 a_in gnd pulse 0 1.8 0 0.1n 0.1n 5n 10n 
v2 b_in gnd pulse 0 1.8 0 0.1n 0.1n 5n 10n 

.tran 0.1n 40n

* Control Statements 
.control
run
plot v(a_in) v(b_in) v(and_out)
print allv > plot_data_v.txt
print alli > plot_data_i.txt
.endc
.end
