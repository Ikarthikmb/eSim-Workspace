* /home/drako/eSim-Workspace/halfadder1/halfadder1.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Jun 29 15:42:13 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  /a /b /sum /carry PORT		
X1  /a /b /carry and_gate		
x1  /a /b /sum xor_gate		

.end
