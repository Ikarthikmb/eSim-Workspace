* /home/drako/esim-workspace/wallace2tree/wallace2tree.cir


.include halfadder.sub
.include and_gate.sub

* u1  a0 a1 b0 b1 z0 z1 z2 z3 port
x1 net-_x1-pad1_ net-_x1-pad2_ z1 net-_x1-pad4_ halfadder
x2 net-_x1-pad4_ net-_x2-pad2_ z2 z3 halfadder
x4 b0 a1 net-_x1-pad2_ and_gate
x3 b0 a0 z0 and_gate
x5 b1 a0 net-_x1-pad1_ and_gate
x6 b1 a1 net-_x2-pad2_ and_gate

v6 b0 0 pulse(0 1.8 0 0.1n 0.1n 5n 10n) 
v3 b1 0 pulse(0 1.8 0 0.1n 0.1n 10n 20n) 
v4 a0 0 pulse(0 1.8 0 0.1n 0.1n 20n 40n)
v5 a1 0 pulse(0 1.8 0 0.1n 0.1n 40n 80n)

.tran 0.1n 80n

* Control Statements 
.control
run
print allv > plot_data_v.txt
print alli > plot_data_i.txt
.endc
.end
