* /home/drako/eSim-Workspace/wallace2tree/wallace2tree.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Jun 29 17:08:21 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  /b0 /a0 /z0 and_gate		
X2  /b0 /a1 Net-_X2-Pad3_ and_gate		
X3  /b1 /a0 Net-_X3-Pad3_ and_gate		
x1  Net-_X3-Pad3_ Net-_X2-Pad3_ /z1 Net-_x1-Pad4_ halfadder		
X4  /b1 /a1 Net-_X4-Pad3_ and_gate		
x2  Net-_x1-Pad4_ Net-_X4-Pad3_ /z2 /z3 halfadder		
U1  /a0 /a1 /b0 /b1 /z0 /z1 /z2 /z3 PORT		

.end
