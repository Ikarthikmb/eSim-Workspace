* /home/drako/applications/eSim-2.1/library/SubcircuitLibrary/halfadder/halfadder.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Jun 29 16:38:50 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ PORT		
X1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad4_ and_gate		
x1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ xor_gate		

.end
