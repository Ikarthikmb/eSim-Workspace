* /home/drako/applications/eSim-2.1/library/SubcircuitLibrary/and_gate/and_gate.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon Jun 28 18:53:16 2021

.lib "~/eSim-Workspace/prelayout/sky130_fd_pr/models/sky130.lib.spice" tt

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M2  Net-_M1-Pad3_ a Net-_M2-Pad3_ Net-_M2-Pad3_ sky130_fd_pr__nfet_01v8 w=1 l=0.5 m=1		
M3  Net-_M2-Pad3_ b GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.5 m=1		
M1  vdd a Net-_M1-Pad3_ vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5 m=1		
M4  vdd b Net-_M1-Pad3_ vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5 m=1		
M5  out Net-_M1-Pad3_ GND GND sky130_fd_pr__nfet_01v8 w=1 l=0.5 m=1		
M6  vdd Net-_M1-Pad3_ out vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5 m=1		
U1  a b out PORT		
v1  vdd GND DC		

.end
